library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.common.all;

entity Nanoprocessor is
    -- port();
end Nanoprocessor;

architecture Behavioral of Nanoprocessor is
begin

end Behavioral;
