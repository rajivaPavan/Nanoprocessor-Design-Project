library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.Logic_Components.Add_Sub_4_bit;

entity AU is
        Port();
end AU;

architecture Behavioral of Add_Sub_4_bit is

begin
    

end Behavioral;

